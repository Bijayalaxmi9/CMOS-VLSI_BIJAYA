***** Spice Netlist for Cell 'Lab9_inverter' *****

************** Module Lab9_inverter **************
.subckt Lab9_inverter vin vout
m1 vout vin gnd gnd scmosn w='0.6u' l='0.4u' m='1' 
m2 vout vin vdd vdd scmosp w='0.6u' l='0.4u' m='1' 
.ends Lab9_inverter




