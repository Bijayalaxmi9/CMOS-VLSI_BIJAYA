***** Spice Netlist for Cell 'Lab9_INV' *****

************** Module Lab9_INV **************
.subckt Lab9_INV vout vin
m2 vout vin vdd vdd scmosp w='0.6u' l='0.4u' m='1' 
m1 vout vin gnd gnd scmosn w='0.6u' l='0.4u' m='1' 
.ends Lab9_INV



